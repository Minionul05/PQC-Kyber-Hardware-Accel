`ifndef DEFINES_VH
`define DEFINES_VH

// CORECT: Spatiu intre nume si valoare. FARA egal, FARA punct si virgula.
`define KYBER_Q 12'd3329
`define DWIDTH 12

`endif